LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY cabine IS 
PORT( 
		E						: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		ET 					: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		AP 					: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		PortOuverte 		: IN STD_LOGIC;
		Horloge 				: IN STD_LOGIC;	
		montee,descend 	: OUT STD_LOGIC; 
		unites,dizaines	: OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
    ); 
END cabine;

ARCHITECTURE ar OF cabine IS

	CONSTANT zero   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000001";
	CONSTANT un     : STD_LOGIC_VECTOR (6 DOWNTO 0) := "1001111";
	CONSTANT deux   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0010010";
	CONSTANT trois  : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000110";
	CONSTANT quatre : STD_LOGIC_VECTOR (6 DOWNTO 0) := "1001100";
	CONSTANT cinq   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0100100";
	CONSTANT six    : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0100000";
	CONSTANT sept   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0001111";
	CONSTANT huit   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000000";
	CONSTANT neuf   : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0000100";
	CONSTANT erreur : STD_LOGIC_VECTOR (6 DOWNTO 0) := "0110000";
	CONSTANT eteint : STD_LOGIC_VECTOR (6 DOWNTO 0) := "1111111";

	TYPE M1_Etat IS (M1_Etat1,M1_Etat2,M1_Etat3,M1_Etat4,M1_Etat5,M1_Etat6,M1_Etat7,M1_Etat8,M1_Etat9,M1_Etat10,M1_Etat11,M1_Etat12,M1_Etat13,M1_Etat14,M1_Etat15,M1_Etat16,M1_Etat17,M1_Etat18,M1_Etat19);
	SIGNAL M1_EtatPresent, M1_EtatSuivant : M1_Etat;

	TYPE M2_Etat IS (M2_Etat1,M2_Etat2,M2_Etat3,M2_Etat4,M2_Etat5);
	SIGNAL M2_EtatPresent, M2_EtatSuivant : M2_Etat;

	SIGNAL ap1Mem : STD_LOGIC;
	SIGNAL ap2Mem : STD_LOGIC;
	SIGNAL ap3Mem : STD_LOGIC;
	SIGNAL ap4Mem : STD_LOGIC;
	SIGNAL finApi : STD_LOGIC;

	BEGIN

	-- DESCRIPTION DU BLOC F
	PROCESS (AP,ET,PortOuverte,ap1Mem,ap2Mem,ap3Mem,ap4Mem)
		BEGIN
		CASE M1_EtatPresent IS
			-- traitement des etages
			WHEN M1_Etat1 => IF ap2Mem='1' OR ap3Mem='1' OR ap4Mem='1' THEN M1_EtatSuivant<=M1_Etat6;
				ELSIF ap1Mem='1' THEN M1_EtatSuivant<=M1_Etat12;
				END IF;
			WHEN M1_Etat2 => IF ap3Mem='1' OR ap4Mem='1' THEN M1_EtatSuivant<=M1_Etat8;
				ELSIF ap2Mem='1' THEN M1_EtatSuivant<=M1_Etat14;
				ELSIF ap1Mem='1' THEN M1_EtatSuivant<=M1_Etat7;
				END IF;
			WHEN M1_Etat3 => IF ap4Mem='1' THEN M1_EtatSuivant<=M1_Etat10;
				ELSIF ap3Mem='1' THEN M1_EtatSuivant<=M1_Etat16;
				ELSIF ap2Mem='1' OR ap1Mem='1' THEN M1_EtatSuivant<=M1_Etat9;
				END IF;
			WHEN M1_Etat4 => IF ap4Mem='1' THEN M1_EtatSuivant<=M1_Etat18;
				ELSIF ap3Mem='1' OR ap2Mem='1' OR ap1Mem='1' THEN M1_EtatSuivant<=M1_Etat11;
				END IF;
				
			--traitement des transistion entre étages
			WHEN M1_Etat5 => IF ET(0)='1' THEN M1_EtatSuivant<=M1_Etat1; END IF;
			WHEN M1_Etat6 => IF ET(1)='1' THEN M1_EtatSuivant<=M1_Etat2; END IF;
			WHEN M1_Etat7 => IF ET(0)='1' THEN M1_EtatSuivant<=M1_Etat1; END IF;
			WHEN M1_Etat8 => IF ET(2)='1' THEN M1_EtatSuivant<=M1_Etat3; END IF;
			WHEN M1_Etat9 => IF ET(1)='1' THEN M1_EtatSuivant<=M1_Etat2; END IF;
			WHEN M1_Etat10 => IF ET(3)='1' THEN M1_EtatSuivant<=M1_Etat4; END IF;
			WHEN M1_Etat11 => IF ET(2)='1' THEN M1_EtatSuivant<=M1_Etat3; END IF;
				
			--traitement des portes
			WHEN M1_Etat12 => IF PortOuverte='1' THEN M1_EtatSuivant<=M1_Etat13; END IF; 	--etage1
			WHEN M1_Etat13 => IF PortOuverte='0' THEN M1_EtatSuivant<=M1_Etat1; END IF; 	--etage1
			WHEN M1_Etat14 => IF PortOuverte='1' THEN M1_EtatSuivant<=M1_Etat15; END IF; 	--etage2
			WHEN M1_Etat15 => IF PortOuverte='0' THEN M1_EtatSuivant<=M1_Etat2; END IF; 	--etage2
			WHEN M1_Etat16 => IF PortOuverte='1' THEN M1_EtatSuivant<=M1_Etat17; END IF; 	--etage3
			WHEN M1_Etat17 => IF PortOuverte='0' THEN M1_EtatSuivant<=M1_Etat3; END IF; 	--etage3
			WHEN M1_Etat18 => IF PortOuverte='1' THEN M1_EtatSuivant<=M1_Etat19; END IF; 	--etage4
			WHEN M1_Etat19 => IF PortOuverte='0' THEN M1_EtatSuivant<=M1_Etat4; END IF; 	--etage4
		END CASE;  
	END PROCESS;
	

	PROCESS (AP,finApi)
		BEGIN
		CASE M2_EtatPresent IS
			WHEN M2_Etat1 => IF finApi='1' THEN M2_EtatSuivant<=M2_Etat5; END IF;
			WHEN M2_Etat2 => IF finApi='1' THEN M2_EtatSuivant<=M2_Etat5; END IF;
			WHEN M2_Etat3 => IF finApi='1' THEN M2_EtatSuivant<=M2_Etat5; END IF;
			WHEN M2_Etat4 => IF finApi='1' THEN M2_EtatSuivant<=M2_Etat5; END IF;
			WHEN M2_Etat5 => 
IF AP(0)='1' THEN M2_EtatSuivant<=M2_Etat1;
				ELSIF AP(1)='1' THEN M2_EtatSuivant<=M2_Etat2;
				ELSIF AP(2)='1' THEN M2_EtatSuivant<=M2_Etat3;
				ELSIF AP(3)='1' THEN M2_EtatSuivant<=M2_Etat4;
				END IF;
		END CASE;
	END PROCESS;

	-- DESCRIPTION DU BLOC M
	PROCESS (Horloge,E) 
	 BEGIN
		-- passage à l'etat suivant
		IF ((Horloge'EVENT) AND (Horloge = '1')) THEN 	M1_EtatPresent <= M1_EtatSuivant; 
M2_EtatPresent <= M2_EtatSuivant; 
		END IF;
		
		-- initialisation des etats
		IF (E(0)='1') THEN M1_EtatPresent<=M1_Etat5; M2_EtatPresent<=M2_Etat5; END IF;
		
	END PROCESS; 

	-- DESCRIPTION DU BLOC G
	-- sorties pour pilotage des afficheurs de la carte
	with M1_EtatPresent select
		unites <= 	zero   	WHEN M1_Etat10,
						un			WHEN M1_Etat1 | M1_Etat11,
						deux		WHEN M1_Etat2 | M1_Etat12,
						trois  	WHEN M1_Etat3 | M1_Etat13,
						quatre 	WHEN M1_Etat4 | M1_Etat14,
						cinq 		WHEN M1_Etat5 | M1_Etat15,
						six		WHEN M1_Etat6 | M1_Etat16,
						sept		WHEN M1_Etat7 | M1_Etat17,
						huit		WHEN M1_Etat8 | M1_Etat18,
						neuf		WHEN M1_Etat9 | M1_Etat19,
						erreur	WHEN OTHERS;
	dizaines <= 	eteint 	WHEN (M1_EtatPresent < M1_Etat10) ELSE 
						un 		WHEN (M1_EtatPresent >= M1_Etat10 AND M1_EtatPresent <= M1_Etat19)ELSE 
						erreur;
		
	-- sorties pour pilotage de la cabine
	montee<='1' WHEN (M1_EtatPresent=M1_Etat6 OR M1_EtatPresent=M1_Etat8 OR M1_EtatPresent=M1_Etat10) ELSE '0';
	descend<='1' WHEN (M1_EtatPresent=M1_Etat7 OR M1_EtatPresent=M1_Etat9 OR M1_EtatPresent=M1_Etat11) ELSE '0';
						
	-- sorties pour memorisation des poussoirs
	ap1Mem<='1' WHEN M2_EtatPresent=M2_Etat1	ELSE '0';
	ap2Mem<='1' WHEN M2_EtatPresent=M2_Etat2	ELSE '0';
	ap3Mem<='1' WHEN M2_EtatPresent=M2_Etat3	ELSE '0';
	ap4Mem<='1' WHEN M2_EtatPresent=M2_Etat4	ELSE '0';

	-- sortie pour mettre fin a ala memorisation du bouton poussoir interne
	WITH M1_EtatPresent select
	finApi <=		'1'	WHEN M1_Etat13 | M1_Etat15 | M1_Etat17 | M1_Etat19,
						'0'	WHEN OTHERS;

END ar;
